magic
tech sky130A
magscale 1 2
timestamp 1700586129
<< nwell >>
rect 1066 349509 558846 349830
rect 1066 348421 558846 348987
rect 1066 347333 558846 347899
rect 1066 346245 558846 346811
rect 1066 345157 558846 345723
rect 1066 344069 558846 344635
rect 1066 342981 558846 343547
rect 1066 341893 558846 342459
rect 1066 340805 558846 341371
rect 1066 339717 558846 340283
rect 1066 338629 558846 339195
rect 1066 337541 558846 338107
rect 1066 336453 558846 337019
rect 1066 335365 558846 335931
rect 1066 334277 558846 334843
rect 1066 333189 558846 333755
rect 1066 332101 558846 332667
rect 1066 331013 558846 331579
rect 1066 329925 558846 330491
rect 1066 328837 558846 329403
rect 1066 327749 558846 328315
rect 1066 326661 558846 327227
rect 1066 325573 558846 326139
rect 1066 324485 558846 325051
rect 1066 323397 558846 323963
rect 1066 322309 558846 322875
rect 1066 321221 558846 321787
rect 1066 320133 558846 320699
rect 1066 319045 558846 319611
rect 1066 317957 558846 318523
rect 1066 316869 558846 317435
rect 1066 315781 558846 316347
rect 1066 314693 558846 315259
rect 1066 313605 558846 314171
rect 1066 312517 558846 313083
rect 1066 311429 558846 311995
rect 1066 310341 558846 310907
rect 1066 309253 558846 309819
rect 1066 308165 558846 308731
rect 1066 307077 558846 307643
rect 1066 305989 558846 306555
rect 1066 304901 558846 305467
rect 1066 303813 558846 304379
rect 1066 302725 558846 303291
rect 1066 301637 558846 302203
rect 1066 300549 558846 301115
rect 1066 299461 558846 300027
rect 1066 298373 558846 298939
rect 1066 297285 558846 297851
rect 1066 296197 558846 296763
rect 1066 295109 558846 295675
rect 1066 294021 558846 294587
rect 1066 292933 558846 293499
rect 1066 291845 558846 292411
rect 1066 290757 558846 291323
rect 1066 289669 558846 290235
rect 1066 288581 558846 289147
rect 1066 287493 558846 288059
rect 1066 286405 558846 286971
rect 1066 285317 558846 285883
rect 1066 284229 558846 284795
rect 1066 283141 558846 283707
rect 1066 282053 558846 282619
rect 1066 280965 558846 281531
rect 1066 279877 558846 280443
rect 1066 278789 558846 279355
rect 1066 277701 558846 278267
rect 1066 276613 558846 277179
rect 1066 275525 558846 276091
rect 1066 274437 558846 275003
rect 1066 273349 558846 273915
rect 1066 272261 558846 272827
rect 1066 271173 558846 271739
rect 1066 270085 558846 270651
rect 1066 268997 558846 269563
rect 1066 267909 558846 268475
rect 1066 266821 558846 267387
rect 1066 265733 558846 266299
rect 1066 264645 558846 265211
rect 1066 263557 558846 264123
rect 1066 262469 558846 263035
rect 1066 261381 558846 261947
rect 1066 260293 558846 260859
rect 1066 259205 558846 259771
rect 1066 258117 558846 258683
rect 1066 257029 558846 257595
rect 1066 255941 558846 256507
rect 1066 254853 558846 255419
rect 1066 253765 558846 254331
rect 1066 252677 558846 253243
rect 1066 251589 558846 252155
rect 1066 250501 558846 251067
rect 1066 249413 558846 249979
rect 1066 248325 558846 248891
rect 1066 247237 558846 247803
rect 1066 246149 558846 246715
rect 1066 245061 558846 245627
rect 1066 243973 558846 244539
rect 1066 242885 558846 243451
rect 1066 241797 558846 242363
rect 1066 240709 558846 241275
rect 1066 239621 558846 240187
rect 1066 238533 558846 239099
rect 1066 237445 558846 238011
rect 1066 236357 558846 236923
rect 1066 235269 558846 235835
rect 1066 234181 558846 234747
rect 1066 233093 558846 233659
rect 1066 232005 558846 232571
rect 1066 230917 558846 231483
rect 1066 229829 558846 230395
rect 1066 228741 558846 229307
rect 1066 227653 558846 228219
rect 1066 226565 558846 227131
rect 1066 225477 558846 226043
rect 1066 224389 558846 224955
rect 1066 223301 558846 223867
rect 1066 222213 558846 222779
rect 1066 221125 558846 221691
rect 1066 220037 558846 220603
rect 1066 218949 558846 219515
rect 1066 217861 558846 218427
rect 1066 216773 558846 217339
rect 1066 215685 558846 216251
rect 1066 214597 558846 215163
rect 1066 213509 558846 214075
rect 1066 212421 558846 212987
rect 1066 211333 558846 211899
rect 1066 210245 558846 210811
rect 1066 209157 558846 209723
rect 1066 208069 558846 208635
rect 1066 206981 558846 207547
rect 1066 205893 558846 206459
rect 1066 204805 558846 205371
rect 1066 203717 558846 204283
rect 1066 202629 558846 203195
rect 1066 201541 558846 202107
rect 1066 200453 558846 201019
rect 1066 199365 558846 199931
rect 1066 198277 558846 198843
rect 1066 197189 558846 197755
rect 1066 196101 558846 196667
rect 1066 195013 558846 195579
rect 1066 193925 558846 194491
rect 1066 192837 558846 193403
rect 1066 191749 558846 192315
rect 1066 190661 558846 191227
rect 1066 189573 558846 190139
rect 1066 188485 558846 189051
rect 1066 187397 558846 187963
rect 1066 186309 558846 186875
rect 1066 185221 558846 185787
rect 1066 184133 558846 184699
rect 1066 183045 558846 183611
rect 1066 181957 558846 182523
rect 1066 180869 558846 181435
rect 1066 179781 558846 180347
rect 1066 178693 558846 179259
rect 1066 177605 558846 178171
rect 1066 176517 558846 177083
rect 1066 175429 558846 175995
rect 1066 174341 558846 174907
rect 1066 173253 558846 173819
rect 1066 172165 558846 172731
rect 1066 171077 558846 171643
rect 1066 169989 558846 170555
rect 1066 168901 558846 169467
rect 1066 167813 558846 168379
rect 1066 166725 558846 167291
rect 1066 165637 558846 166203
rect 1066 164549 558846 165115
rect 1066 163461 558846 164027
rect 1066 162373 558846 162939
rect 1066 161285 558846 161851
rect 1066 160197 558846 160763
rect 1066 159109 558846 159675
rect 1066 158021 558846 158587
rect 1066 156933 558846 157499
rect 1066 155845 558846 156411
rect 1066 154757 558846 155323
rect 1066 153669 558846 154235
rect 1066 152581 558846 153147
rect 1066 151493 558846 152059
rect 1066 150405 558846 150971
rect 1066 149317 558846 149883
rect 1066 148229 558846 148795
rect 1066 147141 558846 147707
rect 1066 146053 558846 146619
rect 1066 144965 558846 145531
rect 1066 143877 558846 144443
rect 1066 142789 558846 143355
rect 1066 141701 558846 142267
rect 1066 140613 558846 141179
rect 1066 139525 558846 140091
rect 1066 138437 558846 139003
rect 1066 137349 558846 137915
rect 1066 136261 558846 136827
rect 1066 135173 558846 135739
rect 1066 134085 558846 134651
rect 1066 132997 558846 133563
rect 1066 131909 558846 132475
rect 1066 130821 558846 131387
rect 1066 129733 558846 130299
rect 1066 128645 558846 129211
rect 1066 127557 558846 128123
rect 1066 126469 558846 127035
rect 1066 125381 558846 125947
rect 1066 124293 558846 124859
rect 1066 123205 558846 123771
rect 1066 122117 558846 122683
rect 1066 121029 558846 121595
rect 1066 119941 558846 120507
rect 1066 118853 558846 119419
rect 1066 117765 558846 118331
rect 1066 116677 558846 117243
rect 1066 115589 558846 116155
rect 1066 114501 558846 115067
rect 1066 113413 558846 113979
rect 1066 112325 558846 112891
rect 1066 111237 558846 111803
rect 1066 110149 558846 110715
rect 1066 109061 558846 109627
rect 1066 107973 558846 108539
rect 1066 106885 558846 107451
rect 1066 105797 558846 106363
rect 1066 104709 558846 105275
rect 1066 103621 558846 104187
rect 1066 102533 558846 103099
rect 1066 101445 558846 102011
rect 1066 100357 558846 100923
rect 1066 99269 558846 99835
rect 1066 98181 558846 98747
rect 1066 97093 558846 97659
rect 1066 96005 558846 96571
rect 1066 94917 558846 95483
rect 1066 93829 558846 94395
rect 1066 92741 558846 93307
rect 1066 91653 558846 92219
rect 1066 90565 558846 91131
rect 1066 89477 558846 90043
rect 1066 88389 558846 88955
rect 1066 87301 558846 87867
rect 1066 86213 558846 86779
rect 1066 85125 558846 85691
rect 1066 84037 558846 84603
rect 1066 82949 558846 83515
rect 1066 81861 558846 82427
rect 1066 80773 558846 81339
rect 1066 79685 558846 80251
rect 1066 78597 558846 79163
rect 1066 77509 558846 78075
rect 1066 76421 558846 76987
rect 1066 75333 558846 75899
rect 1066 74245 558846 74811
rect 1066 73157 558846 73723
rect 1066 72069 558846 72635
rect 1066 70981 558846 71547
rect 1066 69893 558846 70459
rect 1066 68805 558846 69371
rect 1066 67717 558846 68283
rect 1066 66629 558846 67195
rect 1066 65541 558846 66107
rect 1066 64453 558846 65019
rect 1066 63365 558846 63931
rect 1066 62277 558846 62843
rect 1066 61189 558846 61755
rect 1066 60101 558846 60667
rect 1066 59013 558846 59579
rect 1066 57925 558846 58491
rect 1066 56837 558846 57403
rect 1066 55749 558846 56315
rect 1066 54661 558846 55227
rect 1066 53573 558846 54139
rect 1066 52485 558846 53051
rect 1066 51397 558846 51963
rect 1066 50309 558846 50875
rect 1066 49221 558846 49787
rect 1066 48133 558846 48699
rect 1066 47045 558846 47611
rect 1066 45957 558846 46523
rect 1066 44869 558846 45435
rect 1066 43781 558846 44347
rect 1066 42693 558846 43259
rect 1066 41605 558846 42171
rect 1066 40517 558846 41083
rect 1066 39429 558846 39995
rect 1066 38341 558846 38907
rect 1066 37253 558846 37819
rect 1066 36165 558846 36731
rect 1066 35077 558846 35643
rect 1066 33989 558846 34555
rect 1066 32901 558846 33467
rect 1066 31813 558846 32379
rect 1066 30725 558846 31291
rect 1066 29637 558846 30203
rect 1066 28549 558846 29115
rect 1066 27461 558846 28027
rect 1066 26373 558846 26939
rect 1066 25285 558846 25851
rect 1066 24197 558846 24763
rect 1066 23109 558846 23675
rect 1066 22021 558846 22587
rect 1066 20933 558846 21499
rect 1066 19845 558846 20411
rect 1066 18757 558846 19323
rect 1066 17669 558846 18235
rect 1066 16581 558846 17147
rect 1066 15493 558846 16059
rect 1066 14405 558846 14971
rect 1066 13317 558846 13883
rect 1066 12229 558846 12795
rect 1066 11141 558846 11707
rect 1066 10053 558846 10619
rect 1066 8965 558846 9531
rect 1066 7877 558846 8443
rect 1066 6789 558846 7355
rect 1066 5701 558846 6267
rect 1066 4613 558846 5179
rect 1066 3525 558846 4091
rect 1066 2437 558846 3003
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 1104 2128 558978 349840
<< metal2 >>
rect 279974 0 280030 800
<< obsm2 >>
rect 4214 856 558974 349829
rect 4214 800 279918 856
rect 280086 800 558974 856
<< metal3 >>
rect 559200 342184 560000 342304
rect 559200 328312 560000 328432
rect 559200 314440 560000 314560
rect 559200 300568 560000 300688
rect 559200 286696 560000 286816
rect 559200 272824 560000 272944
rect 559200 258952 560000 259072
rect 559200 245080 560000 245200
rect 559200 231208 560000 231328
rect 559200 217336 560000 217456
rect 559200 203464 560000 203584
rect 559200 189592 560000 189712
rect 559200 175720 560000 175840
rect 559200 161848 560000 161968
rect 559200 147976 560000 148096
rect 559200 134104 560000 134224
rect 559200 120232 560000 120352
rect 559200 106360 560000 106480
rect 559200 92488 560000 92608
rect 559200 78616 560000 78736
rect 559200 64744 560000 64864
rect 559200 50872 560000 50992
rect 559200 37000 560000 37120
rect 559200 23128 560000 23248
rect 559200 9256 560000 9376
<< obsm3 >>
rect 4210 342384 559200 349825
rect 4210 342104 559120 342384
rect 4210 328512 559200 342104
rect 4210 328232 559120 328512
rect 4210 314640 559200 328232
rect 4210 314360 559120 314640
rect 4210 300768 559200 314360
rect 4210 300488 559120 300768
rect 4210 286896 559200 300488
rect 4210 286616 559120 286896
rect 4210 273024 559200 286616
rect 4210 272744 559120 273024
rect 4210 259152 559200 272744
rect 4210 258872 559120 259152
rect 4210 245280 559200 258872
rect 4210 245000 559120 245280
rect 4210 231408 559200 245000
rect 4210 231128 559120 231408
rect 4210 217536 559200 231128
rect 4210 217256 559120 217536
rect 4210 203664 559200 217256
rect 4210 203384 559120 203664
rect 4210 189792 559200 203384
rect 4210 189512 559120 189792
rect 4210 175920 559200 189512
rect 4210 175640 559120 175920
rect 4210 162048 559200 175640
rect 4210 161768 559120 162048
rect 4210 148176 559200 161768
rect 4210 147896 559120 148176
rect 4210 134304 559200 147896
rect 4210 134024 559120 134304
rect 4210 120432 559200 134024
rect 4210 120152 559120 120432
rect 4210 106560 559200 120152
rect 4210 106280 559120 106560
rect 4210 92688 559200 106280
rect 4210 92408 559120 92688
rect 4210 78816 559200 92408
rect 4210 78536 559120 78816
rect 4210 64944 559200 78536
rect 4210 64664 559120 64944
rect 4210 51072 559200 64664
rect 4210 50792 559120 51072
rect 4210 37200 559200 50792
rect 4210 36920 559120 37200
rect 4210 23328 559200 36920
rect 4210 23048 559120 23328
rect 4210 9456 559200 23048
rect 4210 9176 559120 9456
rect 4210 2143 559200 9176
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< labels >>
rlabel metal3 s 559200 342184 560000 342304 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 559200 134104 560000 134224 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 559200 120232 560000 120352 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 559200 106360 560000 106480 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 559200 92488 560000 92608 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 559200 78616 560000 78736 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 559200 64744 560000 64864 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 559200 50872 560000 50992 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 559200 37000 560000 37120 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 559200 23128 560000 23248 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 559200 9256 560000 9376 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 559200 314440 560000 314560 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 559200 286696 560000 286816 6 io_in[2]
port 13 nsew signal input
rlabel metal3 s 559200 258952 560000 259072 6 io_in[3]
port 14 nsew signal input
rlabel metal3 s 559200 231208 560000 231328 6 io_in[4]
port 15 nsew signal input
rlabel metal3 s 559200 203464 560000 203584 6 io_in[5]
port 16 nsew signal input
rlabel metal3 s 559200 189592 560000 189712 6 io_in[6]
port 17 nsew signal input
rlabel metal3 s 559200 175720 560000 175840 6 io_in[7]
port 18 nsew signal input
rlabel metal3 s 559200 161848 560000 161968 6 io_in[8]
port 19 nsew signal input
rlabel metal3 s 559200 147976 560000 148096 6 io_in[9]
port 20 nsew signal input
rlabel metal3 s 559200 328312 560000 328432 6 io_out[0]
port 21 nsew signal output
rlabel metal3 s 559200 300568 560000 300688 6 io_out[1]
port 22 nsew signal output
rlabel metal3 s 559200 272824 560000 272944 6 io_out[2]
port 23 nsew signal output
rlabel metal3 s 559200 245080 560000 245200 6 io_out[3]
port 24 nsew signal output
rlabel metal3 s 559200 217336 560000 217456 6 io_out[4]
port 25 nsew signal output
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 26 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 27 nsew ground bidirectional
rlabel metal2 s 279974 0 280030 800 6 wb_clk_i
port 28 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 51690636
string GDS_FILE /home/kiran/special_topic_asics/riscv_control_unit_tapeout/openlane/user_proj_example/runs/23_11_21_22_16/results/signoff/user_proj_example.magic.gds
string GDS_START 199992
<< end >>

