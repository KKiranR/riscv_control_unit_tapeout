VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1710.920 2800.000 1711.520 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 670.520 2800.000 671.120 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 601.160 2800.000 601.760 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 531.800 2800.000 532.400 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 462.440 2800.000 463.040 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 393.080 2800.000 393.680 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 323.720 2800.000 324.320 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 254.360 2800.000 254.960 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 185.000 2800.000 185.600 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 115.640 2800.000 116.240 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 46.280 2800.000 46.880 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1572.200 2800.000 1572.800 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1433.480 2800.000 1434.080 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1294.760 2800.000 1295.360 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1156.040 2800.000 1156.640 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1017.320 2800.000 1017.920 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 947.960 2800.000 948.560 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 878.600 2800.000 879.200 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 809.240 2800.000 809.840 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 739.880 2800.000 740.480 ;
    END
  END io_in[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1641.560 2800.000 1642.160 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1502.840 2800.000 1503.440 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1364.120 2800.000 1364.720 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1225.400 2800.000 1226.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1086.680 2800.000 1087.280 ;
    END
  END io_out[4]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 1749.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 1749.200 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 1399.870 0.000 1400.150 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER nwell ;
        RECT 5.330 1747.545 2794.230 1749.150 ;
        RECT 5.330 1742.105 2794.230 1744.935 ;
        RECT 5.330 1736.665 2794.230 1739.495 ;
        RECT 5.330 1731.225 2794.230 1734.055 ;
        RECT 5.330 1725.785 2794.230 1728.615 ;
        RECT 5.330 1720.345 2794.230 1723.175 ;
        RECT 5.330 1714.905 2794.230 1717.735 ;
        RECT 5.330 1709.465 2794.230 1712.295 ;
        RECT 5.330 1704.025 2794.230 1706.855 ;
        RECT 5.330 1698.585 2794.230 1701.415 ;
        RECT 5.330 1693.145 2794.230 1695.975 ;
        RECT 5.330 1687.705 2794.230 1690.535 ;
        RECT 5.330 1682.265 2794.230 1685.095 ;
        RECT 5.330 1676.825 2794.230 1679.655 ;
        RECT 5.330 1671.385 2794.230 1674.215 ;
        RECT 5.330 1665.945 2794.230 1668.775 ;
        RECT 5.330 1660.505 2794.230 1663.335 ;
        RECT 5.330 1655.065 2794.230 1657.895 ;
        RECT 5.330 1649.625 2794.230 1652.455 ;
        RECT 5.330 1644.185 2794.230 1647.015 ;
        RECT 5.330 1638.745 2794.230 1641.575 ;
        RECT 5.330 1633.305 2794.230 1636.135 ;
        RECT 5.330 1627.865 2794.230 1630.695 ;
        RECT 5.330 1622.425 2794.230 1625.255 ;
        RECT 5.330 1616.985 2794.230 1619.815 ;
        RECT 5.330 1611.545 2794.230 1614.375 ;
        RECT 5.330 1606.105 2794.230 1608.935 ;
        RECT 5.330 1600.665 2794.230 1603.495 ;
        RECT 5.330 1595.225 2794.230 1598.055 ;
        RECT 5.330 1589.785 2794.230 1592.615 ;
        RECT 5.330 1584.345 2794.230 1587.175 ;
        RECT 5.330 1578.905 2794.230 1581.735 ;
        RECT 5.330 1573.465 2794.230 1576.295 ;
        RECT 5.330 1568.025 2794.230 1570.855 ;
        RECT 5.330 1562.585 2794.230 1565.415 ;
        RECT 5.330 1557.145 2794.230 1559.975 ;
        RECT 5.330 1551.705 2794.230 1554.535 ;
        RECT 5.330 1546.265 2794.230 1549.095 ;
        RECT 5.330 1540.825 2794.230 1543.655 ;
        RECT 5.330 1535.385 2794.230 1538.215 ;
        RECT 5.330 1529.945 2794.230 1532.775 ;
        RECT 5.330 1524.505 2794.230 1527.335 ;
        RECT 5.330 1519.065 2794.230 1521.895 ;
        RECT 5.330 1513.625 2794.230 1516.455 ;
        RECT 5.330 1508.185 2794.230 1511.015 ;
        RECT 5.330 1502.745 2794.230 1505.575 ;
        RECT 5.330 1497.305 2794.230 1500.135 ;
        RECT 5.330 1491.865 2794.230 1494.695 ;
        RECT 5.330 1486.425 2794.230 1489.255 ;
        RECT 5.330 1480.985 2794.230 1483.815 ;
        RECT 5.330 1475.545 2794.230 1478.375 ;
        RECT 5.330 1470.105 2794.230 1472.935 ;
        RECT 5.330 1464.665 2794.230 1467.495 ;
        RECT 5.330 1459.225 2794.230 1462.055 ;
        RECT 5.330 1453.785 2794.230 1456.615 ;
        RECT 5.330 1448.345 2794.230 1451.175 ;
        RECT 5.330 1442.905 2794.230 1445.735 ;
        RECT 5.330 1437.465 2794.230 1440.295 ;
        RECT 5.330 1432.025 2794.230 1434.855 ;
        RECT 5.330 1426.585 2794.230 1429.415 ;
        RECT 5.330 1421.145 2794.230 1423.975 ;
        RECT 5.330 1415.705 2794.230 1418.535 ;
        RECT 5.330 1410.265 2794.230 1413.095 ;
        RECT 5.330 1404.825 2794.230 1407.655 ;
        RECT 5.330 1399.385 2794.230 1402.215 ;
        RECT 5.330 1393.945 2794.230 1396.775 ;
        RECT 5.330 1388.505 2794.230 1391.335 ;
        RECT 5.330 1383.065 2794.230 1385.895 ;
        RECT 5.330 1377.625 2794.230 1380.455 ;
        RECT 5.330 1372.185 2794.230 1375.015 ;
        RECT 5.330 1366.745 2794.230 1369.575 ;
        RECT 5.330 1361.305 2794.230 1364.135 ;
        RECT 5.330 1355.865 2794.230 1358.695 ;
        RECT 5.330 1350.425 2794.230 1353.255 ;
        RECT 5.330 1344.985 2794.230 1347.815 ;
        RECT 5.330 1339.545 2794.230 1342.375 ;
        RECT 5.330 1334.105 2794.230 1336.935 ;
        RECT 5.330 1328.665 2794.230 1331.495 ;
        RECT 5.330 1323.225 2794.230 1326.055 ;
        RECT 5.330 1317.785 2794.230 1320.615 ;
        RECT 5.330 1312.345 2794.230 1315.175 ;
        RECT 5.330 1306.905 2794.230 1309.735 ;
        RECT 5.330 1301.465 2794.230 1304.295 ;
        RECT 5.330 1296.025 2794.230 1298.855 ;
        RECT 5.330 1290.585 2794.230 1293.415 ;
        RECT 5.330 1285.145 2794.230 1287.975 ;
        RECT 5.330 1279.705 2794.230 1282.535 ;
        RECT 5.330 1274.265 2794.230 1277.095 ;
        RECT 5.330 1268.825 2794.230 1271.655 ;
        RECT 5.330 1263.385 2794.230 1266.215 ;
        RECT 5.330 1257.945 2794.230 1260.775 ;
        RECT 5.330 1252.505 2794.230 1255.335 ;
        RECT 5.330 1247.065 2794.230 1249.895 ;
        RECT 5.330 1241.625 2794.230 1244.455 ;
        RECT 5.330 1236.185 2794.230 1239.015 ;
        RECT 5.330 1230.745 2794.230 1233.575 ;
        RECT 5.330 1225.305 2794.230 1228.135 ;
        RECT 5.330 1219.865 2794.230 1222.695 ;
        RECT 5.330 1214.425 2794.230 1217.255 ;
        RECT 5.330 1208.985 2794.230 1211.815 ;
        RECT 5.330 1203.545 2794.230 1206.375 ;
        RECT 5.330 1198.105 2794.230 1200.935 ;
        RECT 5.330 1192.665 2794.230 1195.495 ;
        RECT 5.330 1187.225 2794.230 1190.055 ;
        RECT 5.330 1181.785 2794.230 1184.615 ;
        RECT 5.330 1176.345 2794.230 1179.175 ;
        RECT 5.330 1170.905 2794.230 1173.735 ;
        RECT 5.330 1165.465 2794.230 1168.295 ;
        RECT 5.330 1160.025 2794.230 1162.855 ;
        RECT 5.330 1154.585 2794.230 1157.415 ;
        RECT 5.330 1149.145 2794.230 1151.975 ;
        RECT 5.330 1143.705 2794.230 1146.535 ;
        RECT 5.330 1138.265 2794.230 1141.095 ;
        RECT 5.330 1132.825 2794.230 1135.655 ;
        RECT 5.330 1127.385 2794.230 1130.215 ;
        RECT 5.330 1121.945 2794.230 1124.775 ;
        RECT 5.330 1116.505 2794.230 1119.335 ;
        RECT 5.330 1111.065 2794.230 1113.895 ;
        RECT 5.330 1105.625 2794.230 1108.455 ;
        RECT 5.330 1100.185 2794.230 1103.015 ;
        RECT 5.330 1094.745 2794.230 1097.575 ;
        RECT 5.330 1089.305 2794.230 1092.135 ;
        RECT 5.330 1083.865 2794.230 1086.695 ;
        RECT 5.330 1078.425 2794.230 1081.255 ;
        RECT 5.330 1072.985 2794.230 1075.815 ;
        RECT 5.330 1067.545 2794.230 1070.375 ;
        RECT 5.330 1062.105 2794.230 1064.935 ;
        RECT 5.330 1056.665 2794.230 1059.495 ;
        RECT 5.330 1051.225 2794.230 1054.055 ;
        RECT 5.330 1045.785 2794.230 1048.615 ;
        RECT 5.330 1040.345 2794.230 1043.175 ;
        RECT 5.330 1034.905 2794.230 1037.735 ;
        RECT 5.330 1029.465 2794.230 1032.295 ;
        RECT 5.330 1024.025 2794.230 1026.855 ;
        RECT 5.330 1018.585 2794.230 1021.415 ;
        RECT 5.330 1013.145 2794.230 1015.975 ;
        RECT 5.330 1007.705 2794.230 1010.535 ;
        RECT 5.330 1002.265 2794.230 1005.095 ;
        RECT 5.330 996.825 2794.230 999.655 ;
        RECT 5.330 991.385 2794.230 994.215 ;
        RECT 5.330 985.945 2794.230 988.775 ;
        RECT 5.330 980.505 2794.230 983.335 ;
        RECT 5.330 975.065 2794.230 977.895 ;
        RECT 5.330 969.625 2794.230 972.455 ;
        RECT 5.330 964.185 2794.230 967.015 ;
        RECT 5.330 958.745 2794.230 961.575 ;
        RECT 5.330 953.305 2794.230 956.135 ;
        RECT 5.330 947.865 2794.230 950.695 ;
        RECT 5.330 942.425 2794.230 945.255 ;
        RECT 5.330 936.985 2794.230 939.815 ;
        RECT 5.330 931.545 2794.230 934.375 ;
        RECT 5.330 926.105 2794.230 928.935 ;
        RECT 5.330 920.665 2794.230 923.495 ;
        RECT 5.330 915.225 2794.230 918.055 ;
        RECT 5.330 909.785 2794.230 912.615 ;
        RECT 5.330 904.345 2794.230 907.175 ;
        RECT 5.330 898.905 2794.230 901.735 ;
        RECT 5.330 893.465 2794.230 896.295 ;
        RECT 5.330 888.025 2794.230 890.855 ;
        RECT 5.330 882.585 2794.230 885.415 ;
        RECT 5.330 877.145 2794.230 879.975 ;
        RECT 5.330 871.705 2794.230 874.535 ;
        RECT 5.330 866.265 2794.230 869.095 ;
        RECT 5.330 860.825 2794.230 863.655 ;
        RECT 5.330 855.385 2794.230 858.215 ;
        RECT 5.330 849.945 2794.230 852.775 ;
        RECT 5.330 844.505 2794.230 847.335 ;
        RECT 5.330 839.065 2794.230 841.895 ;
        RECT 5.330 833.625 2794.230 836.455 ;
        RECT 5.330 828.185 2794.230 831.015 ;
        RECT 5.330 822.745 2794.230 825.575 ;
        RECT 5.330 817.305 2794.230 820.135 ;
        RECT 5.330 811.865 2794.230 814.695 ;
        RECT 5.330 806.425 2794.230 809.255 ;
        RECT 5.330 800.985 2794.230 803.815 ;
        RECT 5.330 795.545 2794.230 798.375 ;
        RECT 5.330 790.105 2794.230 792.935 ;
        RECT 5.330 784.665 2794.230 787.495 ;
        RECT 5.330 779.225 2794.230 782.055 ;
        RECT 5.330 773.785 2794.230 776.615 ;
        RECT 5.330 768.345 2794.230 771.175 ;
        RECT 5.330 762.905 2794.230 765.735 ;
        RECT 5.330 757.465 2794.230 760.295 ;
        RECT 5.330 752.025 2794.230 754.855 ;
        RECT 5.330 746.585 2794.230 749.415 ;
        RECT 5.330 741.145 2794.230 743.975 ;
        RECT 5.330 735.705 2794.230 738.535 ;
        RECT 5.330 730.265 2794.230 733.095 ;
        RECT 5.330 724.825 2794.230 727.655 ;
        RECT 5.330 719.385 2794.230 722.215 ;
        RECT 5.330 713.945 2794.230 716.775 ;
        RECT 5.330 708.505 2794.230 711.335 ;
        RECT 5.330 703.065 2794.230 705.895 ;
        RECT 5.330 697.625 2794.230 700.455 ;
        RECT 5.330 692.185 2794.230 695.015 ;
        RECT 5.330 686.745 2794.230 689.575 ;
        RECT 5.330 681.305 2794.230 684.135 ;
        RECT 5.330 675.865 2794.230 678.695 ;
        RECT 5.330 670.425 2794.230 673.255 ;
        RECT 5.330 664.985 2794.230 667.815 ;
        RECT 5.330 659.545 2794.230 662.375 ;
        RECT 5.330 654.105 2794.230 656.935 ;
        RECT 5.330 648.665 2794.230 651.495 ;
        RECT 5.330 643.225 2794.230 646.055 ;
        RECT 5.330 637.785 2794.230 640.615 ;
        RECT 5.330 632.345 2794.230 635.175 ;
        RECT 5.330 626.905 2794.230 629.735 ;
        RECT 5.330 621.465 2794.230 624.295 ;
        RECT 5.330 616.025 2794.230 618.855 ;
        RECT 5.330 610.585 2794.230 613.415 ;
        RECT 5.330 605.145 2794.230 607.975 ;
        RECT 5.330 599.705 2794.230 602.535 ;
        RECT 5.330 594.265 2794.230 597.095 ;
        RECT 5.330 588.825 2794.230 591.655 ;
        RECT 5.330 583.385 2794.230 586.215 ;
        RECT 5.330 577.945 2794.230 580.775 ;
        RECT 5.330 572.505 2794.230 575.335 ;
        RECT 5.330 567.065 2794.230 569.895 ;
        RECT 5.330 561.625 2794.230 564.455 ;
        RECT 5.330 556.185 2794.230 559.015 ;
        RECT 5.330 550.745 2794.230 553.575 ;
        RECT 5.330 545.305 2794.230 548.135 ;
        RECT 5.330 539.865 2794.230 542.695 ;
        RECT 5.330 534.425 2794.230 537.255 ;
        RECT 5.330 528.985 2794.230 531.815 ;
        RECT 5.330 523.545 2794.230 526.375 ;
        RECT 5.330 518.105 2794.230 520.935 ;
        RECT 5.330 512.665 2794.230 515.495 ;
        RECT 5.330 507.225 2794.230 510.055 ;
        RECT 5.330 501.785 2794.230 504.615 ;
        RECT 5.330 496.345 2794.230 499.175 ;
        RECT 5.330 490.905 2794.230 493.735 ;
        RECT 5.330 485.465 2794.230 488.295 ;
        RECT 5.330 480.025 2794.230 482.855 ;
        RECT 5.330 474.585 2794.230 477.415 ;
        RECT 5.330 469.145 2794.230 471.975 ;
        RECT 5.330 463.705 2794.230 466.535 ;
        RECT 5.330 458.265 2794.230 461.095 ;
        RECT 5.330 452.825 2794.230 455.655 ;
        RECT 5.330 447.385 2794.230 450.215 ;
        RECT 5.330 441.945 2794.230 444.775 ;
        RECT 5.330 436.505 2794.230 439.335 ;
        RECT 5.330 431.065 2794.230 433.895 ;
        RECT 5.330 425.625 2794.230 428.455 ;
        RECT 5.330 420.185 2794.230 423.015 ;
        RECT 5.330 414.745 2794.230 417.575 ;
        RECT 5.330 409.305 2794.230 412.135 ;
        RECT 5.330 403.865 2794.230 406.695 ;
        RECT 5.330 398.425 2794.230 401.255 ;
        RECT 5.330 392.985 2794.230 395.815 ;
        RECT 5.330 387.545 2794.230 390.375 ;
        RECT 5.330 382.105 2794.230 384.935 ;
        RECT 5.330 376.665 2794.230 379.495 ;
        RECT 5.330 371.225 2794.230 374.055 ;
        RECT 5.330 365.785 2794.230 368.615 ;
        RECT 5.330 360.345 2794.230 363.175 ;
        RECT 5.330 354.905 2794.230 357.735 ;
        RECT 5.330 349.465 2794.230 352.295 ;
        RECT 5.330 344.025 2794.230 346.855 ;
        RECT 5.330 338.585 2794.230 341.415 ;
        RECT 5.330 333.145 2794.230 335.975 ;
        RECT 5.330 327.705 2794.230 330.535 ;
        RECT 5.330 322.265 2794.230 325.095 ;
        RECT 5.330 316.825 2794.230 319.655 ;
        RECT 5.330 311.385 2794.230 314.215 ;
        RECT 5.330 305.945 2794.230 308.775 ;
        RECT 5.330 300.505 2794.230 303.335 ;
        RECT 5.330 295.065 2794.230 297.895 ;
        RECT 5.330 289.625 2794.230 292.455 ;
        RECT 5.330 284.185 2794.230 287.015 ;
        RECT 5.330 278.745 2794.230 281.575 ;
        RECT 5.330 273.305 2794.230 276.135 ;
        RECT 5.330 267.865 2794.230 270.695 ;
        RECT 5.330 262.425 2794.230 265.255 ;
        RECT 5.330 256.985 2794.230 259.815 ;
        RECT 5.330 251.545 2794.230 254.375 ;
        RECT 5.330 246.105 2794.230 248.935 ;
        RECT 5.330 240.665 2794.230 243.495 ;
        RECT 5.330 235.225 2794.230 238.055 ;
        RECT 5.330 229.785 2794.230 232.615 ;
        RECT 5.330 224.345 2794.230 227.175 ;
        RECT 5.330 218.905 2794.230 221.735 ;
        RECT 5.330 213.465 2794.230 216.295 ;
        RECT 5.330 208.025 2794.230 210.855 ;
        RECT 5.330 202.585 2794.230 205.415 ;
        RECT 5.330 197.145 2794.230 199.975 ;
        RECT 5.330 191.705 2794.230 194.535 ;
        RECT 5.330 186.265 2794.230 189.095 ;
        RECT 5.330 180.825 2794.230 183.655 ;
        RECT 5.330 175.385 2794.230 178.215 ;
        RECT 5.330 169.945 2794.230 172.775 ;
        RECT 5.330 164.505 2794.230 167.335 ;
        RECT 5.330 159.065 2794.230 161.895 ;
        RECT 5.330 153.625 2794.230 156.455 ;
        RECT 5.330 148.185 2794.230 151.015 ;
        RECT 5.330 142.745 2794.230 145.575 ;
        RECT 5.330 137.305 2794.230 140.135 ;
        RECT 5.330 131.865 2794.230 134.695 ;
        RECT 5.330 126.425 2794.230 129.255 ;
        RECT 5.330 120.985 2794.230 123.815 ;
        RECT 5.330 115.545 2794.230 118.375 ;
        RECT 5.330 110.105 2794.230 112.935 ;
        RECT 5.330 104.665 2794.230 107.495 ;
        RECT 5.330 99.225 2794.230 102.055 ;
        RECT 5.330 93.785 2794.230 96.615 ;
        RECT 5.330 88.345 2794.230 91.175 ;
        RECT 5.330 82.905 2794.230 85.735 ;
        RECT 5.330 77.465 2794.230 80.295 ;
        RECT 5.330 72.025 2794.230 74.855 ;
        RECT 5.330 66.585 2794.230 69.415 ;
        RECT 5.330 61.145 2794.230 63.975 ;
        RECT 5.330 55.705 2794.230 58.535 ;
        RECT 5.330 50.265 2794.230 53.095 ;
        RECT 5.330 44.825 2794.230 47.655 ;
        RECT 5.330 39.385 2794.230 42.215 ;
        RECT 5.330 33.945 2794.230 36.775 ;
        RECT 5.330 28.505 2794.230 31.335 ;
        RECT 5.330 23.065 2794.230 25.895 ;
        RECT 5.330 17.625 2794.230 20.455 ;
        RECT 5.330 12.185 2794.230 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 1749.045 ;
      LAYER met1 ;
        RECT 5.520 10.640 2794.890 1749.200 ;
      LAYER met2 ;
        RECT 21.070 4.280 2794.870 1749.145 ;
        RECT 21.070 4.000 1399.590 4.280 ;
        RECT 1400.430 4.000 2794.870 4.280 ;
      LAYER met3 ;
        RECT 21.050 1711.920 2796.000 1749.125 ;
        RECT 21.050 1710.520 2795.600 1711.920 ;
        RECT 21.050 1642.560 2796.000 1710.520 ;
        RECT 21.050 1641.160 2795.600 1642.560 ;
        RECT 21.050 1573.200 2796.000 1641.160 ;
        RECT 21.050 1571.800 2795.600 1573.200 ;
        RECT 21.050 1503.840 2796.000 1571.800 ;
        RECT 21.050 1502.440 2795.600 1503.840 ;
        RECT 21.050 1434.480 2796.000 1502.440 ;
        RECT 21.050 1433.080 2795.600 1434.480 ;
        RECT 21.050 1365.120 2796.000 1433.080 ;
        RECT 21.050 1363.720 2795.600 1365.120 ;
        RECT 21.050 1295.760 2796.000 1363.720 ;
        RECT 21.050 1294.360 2795.600 1295.760 ;
        RECT 21.050 1226.400 2796.000 1294.360 ;
        RECT 21.050 1225.000 2795.600 1226.400 ;
        RECT 21.050 1157.040 2796.000 1225.000 ;
        RECT 21.050 1155.640 2795.600 1157.040 ;
        RECT 21.050 1087.680 2796.000 1155.640 ;
        RECT 21.050 1086.280 2795.600 1087.680 ;
        RECT 21.050 1018.320 2796.000 1086.280 ;
        RECT 21.050 1016.920 2795.600 1018.320 ;
        RECT 21.050 948.960 2796.000 1016.920 ;
        RECT 21.050 947.560 2795.600 948.960 ;
        RECT 21.050 879.600 2796.000 947.560 ;
        RECT 21.050 878.200 2795.600 879.600 ;
        RECT 21.050 810.240 2796.000 878.200 ;
        RECT 21.050 808.840 2795.600 810.240 ;
        RECT 21.050 740.880 2796.000 808.840 ;
        RECT 21.050 739.480 2795.600 740.880 ;
        RECT 21.050 671.520 2796.000 739.480 ;
        RECT 21.050 670.120 2795.600 671.520 ;
        RECT 21.050 602.160 2796.000 670.120 ;
        RECT 21.050 600.760 2795.600 602.160 ;
        RECT 21.050 532.800 2796.000 600.760 ;
        RECT 21.050 531.400 2795.600 532.800 ;
        RECT 21.050 463.440 2796.000 531.400 ;
        RECT 21.050 462.040 2795.600 463.440 ;
        RECT 21.050 394.080 2796.000 462.040 ;
        RECT 21.050 392.680 2795.600 394.080 ;
        RECT 21.050 324.720 2796.000 392.680 ;
        RECT 21.050 323.320 2795.600 324.720 ;
        RECT 21.050 255.360 2796.000 323.320 ;
        RECT 21.050 253.960 2795.600 255.360 ;
        RECT 21.050 186.000 2796.000 253.960 ;
        RECT 21.050 184.600 2795.600 186.000 ;
        RECT 21.050 116.640 2796.000 184.600 ;
        RECT 21.050 115.240 2795.600 116.640 ;
        RECT 21.050 47.280 2796.000 115.240 ;
        RECT 21.050 45.880 2795.600 47.280 ;
        RECT 21.050 10.715 2796.000 45.880 ;
  END
END user_proj_example
END LIBRARY

